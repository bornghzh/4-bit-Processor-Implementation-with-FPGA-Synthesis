
module Zarb(
	input [3:0] A,
	input [3:0] B,
	output [7:0] F
    );
	and(F[0],A[0],B[0]);
	and(w1_1,A[1],B[0]);
	and(w1_2,A[2],B[0]);
	and(w1_3,A[3],B[0]);

	and(w1_4,A[0],B[1]);
	and(w1_5,A[1],B[1]);
	and(w1_6,A[2],B[1]);
	and(w1_7,A[3],B[1]);

FA4 S1 ({1'b0,w1_3,w1_2,w1_1},{w1_7,w1_6,w1_5,w1_4},{g1_4,g1_3,g1_2,g1_1,F[1]});

	and(w2_1,A[0],B[2]);
	and(w2_2,A[1],B[2]);
	and(w2_3,A[2],B[2]);
	and(w2_4,A[3],B[2]);

FA4 S2 ({g1_4,g1_3,g1_2,g1_1},{w2_4,w2_3,w2_2,w2_1},{g2_4,g2_3,g2_2,g2_1,F[2]});
	 
	and(w3_1,A[0],B[3]);
	and(w3_2,A[1],B[3]);
	and(w3_3,A[2],B[3]);
	and(w3_4,A[3],B[3]);

FA4 S3 ({g2_4,g2_3,g2_2,g2_1},{w3_4,w3_3,w3_2,w3_1},{F[7],F[6],F[5],F[4],F[3]});


endmodule
